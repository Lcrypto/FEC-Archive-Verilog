//
// Project       : ccsds turbo
// Author        : Shekhalev Denis (des00)
// Workfile      : ccsds_parameters.vh
// Description   :
//

  localparam int cN_TAB  [4] = '{223*8*1, 223*8*2, 223*8*4, 223*8*5};

  //------------------------------------------------------------------------------------------------------
  // permutation address logic base data width
  //------------------------------------------------------------------------------------------------------

  parameter int cW = 14;  // don't change

  typedef logic [cW-1 : 0] ptab_dat_t;

  //------------------------------------------------------------------------------------------------------
  //
  //------------------------------------------------------------------------------------------------------

  //
  // code constants to use instead of digits
  typedef enum bit [1 : 0] {
    cCODE_1by2  = 2'h0,
    cCODE_1by3  = 2'h1,
    cCODE_1by4  = 2'h2,
    cCODE_1by6  = 2'h3
  } ccsds_turbo_code_t;

  //------------------------------------------------------------------------------------------------------
  //
  //------------------------------------------------------------------------------------------------------
