//
// (!!!) IT'S GENERATED short table for 7/8 coderate, 8176 bits do 1 LLR per cycle(!!!)
//
  addr_tab[0][0][0][0] = '{baddr:0, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][0][1][0] = '{baddr:12, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][0][2][0] = '{baddr:0, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][0][3][0] = '{baddr:24, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][0][4][0] = '{baddr:0, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][0][5][0] = '{baddr:151, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][0][6][0] = '{baddr:0, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][0][7][0] = '{baddr:9, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][0][8][0] = '{baddr:0, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][0][9][0] = '{baddr:53, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][0][10][0] = '{baddr:0, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][0][11][0] = '{baddr:18, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][0][12][0] = '{baddr:0, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][0][13][0] = '{baddr:202, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][0][14][0] = '{baddr:0, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][0][15][0] = '{baddr:36, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][1][0][0] = '{baddr:176, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][1][1][0] = '{baddr:239, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][1][2][0] = '{baddr:352, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][1][3][0] = '{baddr:431, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][1][4][0] = '{baddr:392, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][1][5][0] = '{baddr:409, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][1][6][0] = '{baddr:351, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][1][7][0] = '{baddr:359, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][1][8][0] = '{baddr:307, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][1][9][0] = '{baddr:329, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][1][10][0] = '{baddr:207, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][1][11][0] = '{baddr:281, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][1][12][0] = '{baddr:399, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][1][13][0] = '{baddr:457, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][1][14][0] = '{baddr:247, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[0][1][15][0] = '{baddr:261, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][0][0][0] = '{baddr:99, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][0][1][0] = '{baddr:130, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][0][2][0] = '{baddr:198, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][0][3][0] = '{baddr:260, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][0][4][0] = '{baddr:215, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][0][5][0] = '{baddr:282, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][0][6][0] = '{baddr:48, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][0][7][0] = '{baddr:193, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][0][8][0] = '{baddr:273, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][0][9][0] = '{baddr:302, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][0][10][0] = '{baddr:96, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][0][11][0] = '{baddr:191, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][0][12][0] = '{baddr:244, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][0][13][0] = '{baddr:364, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][0][14][0] = '{baddr:51, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][0][15][0] = '{baddr:192, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][1][0][0] = '{baddr:471, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][1][1][0] = '{baddr:473, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][1][2][0] = '{baddr:435, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][1][3][0] = '{baddr:478, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][1][4][0] = '{baddr:420, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][1][5][0] = '{baddr:481, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][1][6][0] = '{baddr:396, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][1][7][0] = '{baddr:445, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][1][8][0] = '{baddr:430, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][1][9][0] = '{baddr:451, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][1][10][0] = '{baddr:379, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][1][11][0] = '{baddr:386, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][1][12][0] = '{baddr:467, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][1][13][0] = '{baddr:470, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][1][14][0] = '{baddr:382, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
  addr_tab[1][1][15][0] = '{baddr:414, offset:'{0}, offsetm:'{0}, sela:'{0}, invsela:'{0}};
