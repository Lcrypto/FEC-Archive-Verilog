/*






  logic          gaus_log_tab__iclk     ;
  logic          gaus_log_tab__ireset   ;
  logic          gaus_log_tab__iclkena  ;
  logic  [8 : 0] gaus_log_tab__iaddr0   ;
  logic  [8 : 0] gaus_log_tab__iaddr1   ;
  logic [17 : 0] gaus_log_tab__odat0    ;
  logic [17 : 0] gaus_log_tab__odat1    ;



  gaus_log_tab
  gaus_log_tab
  (
    .iclk    ( gaus_log_tab__iclk    ) ,
    .ireset  ( gaus_log_tab__ireset  ) ,
    .iclkena ( gaus_log_tab__iclkena ) ,
    .iaddr0  ( gaus_log_tab__iaddr0  ) ,
    .iaddr1  ( gaus_log_tab__iaddr1  ) ,
    .odat0   ( gaus_log_tab__odat0   ) ,
    .odat1   ( gaus_log_tab__odat1   )
  );


  assign gaus_log_tab__iclk    = '0 ;
  assign gaus_log_tab__ireset  = '0 ;
  assign gaus_log_tab__iclkena = '0 ;
  assign gaus_log_tab__iaddr0  = '0 ;
  assign gaus_log_tab__iaddr1  = '0 ;



*/


//
// Project       : gaus_log_tab
// Author        : Shekhalev Denis (des00)
// Revision      : $Revision$
// Date          : $Date$
// Workfile      : gaus_log_tab.v
// Description   : ROM based sqrt(log) for simple Box-Muller algorithm
//

module gaus_log_tab
(
  iclk    ,
  ireset  ,
  iclkena ,
  //
  iaddr0  ,
  iaddr1  ,
  //
  odat0   ,
  odat1
);

  //------------------------------------------------------------------------------------------------------
  //
  //------------------------------------------------------------------------------------------------------

  input  logic          iclk     ;
  input  logic          ireset   ;
  input  logic          iclkena  ;
  //
  input  logic  [8 : 0] iaddr0   ;
  input  logic  [8 : 0] iaddr1   ;
  //
  output logic [17 : 0] odat0    ;
  output logic [17 : 0] odat1    ;

  //------------------------------------------------------------------------------------------------------
  //
  //------------------------------------------------------------------------------------------------------

  localparam logic signed [17 : 0] cLOG_TAB [0 : 511] = '{
    130950,
    123460,
    118861,
    115487,
    112800,
    110556,
    108623,
    106920,
    105395,
    104012,
    102745,
    101574,
    100485,
    99467,
    98509,
    97604,
    96747,
    95931,
    95153,
    94410,
    93697,
    93012,
    92353,
    91717,
    91103,
    90510,
    89935,
    89377,
    88836,
    88310,
    87798,
    87300,
    86814,
    86340,
    85877,
    85425,
    84983,
    84551,
    84128,
    83713,
    83307,
    82908,
    82517,
    82133,
    81756,
    81386,
    81022,
    80664,
    80312,
    79966,
    79624,
    79289,
    78958,
    78632,
    78310,
    77993,
    77681,
    77373,
    77068,
    76768,
    76472,
    76179,
    75889,
    75604,
    75321,
    75042,
    74766,
    74494,
    74224,
    73957,
    73693,
    73431,
    73173,
    72917,
    72663,
    72412,
    72164,
    71918,
    71674,
    71432,
    71193,
    70955,
    70720,
    70487,
    70256,
    70027,
    69800,
    69574,
    69351,
    69129,
    68909,
    68690,
    68474,
    68259,
    68045,
    67834,
    67623,
    67414,
    67207,
    67001,
    66797,
    66594,
    66392,
    66192,
    65993,
    65795,
    65599,
    65404,
    65210,
    65017,
    64825,
    64635,
    64446,
    64257,
    64070,
    63884,
    63699,
    63515,
    63333,
    63151,
    62970,
    62790,
    62611,
    62433,
    62256,
    62080,
    61905,
    61730,
    61557,
    61384,
    61212,
    61041,
    60871,
    60702,
    60533,
    60365,
    60198,
    60032,
    59866,
    59702,
    59538,
    59374,
    59212,
    59050,
    58888,
    58728,
    58568,
    58408,
    58250,
    58092,
    57934,
    57777,
    57621,
    57466,
    57311,
    57156,
    57002,
    56849,
    56696,
    56544,
    56393,
    56241,
    56091,
    55941,
    55791,
    55642,
    55494,
    55346,
    55198,
    55051,
    54904,
    54758,
    54612,
    54467,
    54322,
    54178,
    54034,
    53891,
    53748,
    53605,
    53463,
    53321,
    53179,
    53038,
    52898,
    52757,
    52618,
    52478,
    52339,
    52200,
    52062,
    51924,
    51786,
    51649,
    51512,
    51375,
    51239,
    51103,
    50967,
    50832,
    50697,
    50562,
    50428,
    50294,
    50160,
    50026,
    49893,
    49760,
    49627,
    49495,
    49363,
    49231,
    49100,
    48968,
    48837,
    48707,
    48576,
    48446,
    48316,
    48186,
    48056,
    47927,
    47798,
    47669,
    47541,
    47412,
    47284,
    47156,
    47028,
    46901,
    46774,
    46647,
    46520,
    46393,
    46266,
    46140,
    46014,
    45888,
    45762,
    45637,
    45511,
    45386,
    45261,
    45136,
    45011,
    44887,
    44763,
    44638,
    44514,
    44390,
    44267,
    44143,
    44019,
    43896,
    43773,
    43650,
    43527,
    43404,
    43281,
    43159,
    43036,
    42914,
    42792,
    42670,
    42548,
    42426,
    42304,
    42183,
    42061,
    41940,
    41819,
    41697,
    41576,
    41455,
    41334,
    41213,
    41093,
    40972,
    40851,
    40731,
    40610,
    40490,
    40369,
    40249,
    40129,
    40009,
    39889,
    39769,
    39649,
    39529,
    39409,
    39289,
    39169,
    39050,
    38930,
    38810,
    38691,
    38571,
    38451,
    38332,
    38212,
    38093,
    37974,
    37854,
    37735,
    37615,
    37496,
    37376,
    37257,
    37138,
    37018,
    36899,
    36780,
    36660,
    36541,
    36421,
    36302,
    36182,
    36063,
    35944,
    35824,
    35704,
    35585,
    35465,
    35346,
    35226,
    35106,
    34987,
    34867,
    34747,
    34627,
    34507,
    34387,
    34267,
    34147,
    34027,
    33907,
    33786,
    33666,
    33545,
    33425,
    33304,
    33184,
    33063,
    32942,
    32821,
    32700,
    32579,
    32457,
    32336,
    32214,
    32093,
    31971,
    31849,
    31727,
    31605,
    31483,
    31361,
    31238,
    31116,
    30993,
    30870,
    30747,
    30624,
    30500,
    30377,
    30253,
    30129,
    30005,
    29881,
    29756,
    29632,
    29507,
    29382,
    29257,
    29132,
    29006,
    28880,
    28754,
    28628,
    28501,
    28375,
    28248,
    28121,
    27993,
    27866,
    27738,
    27610,
    27481,
    27352,
    27223,
    27094,
    26965,
    26835,
    26705,
    26574,
    26443,
    26312,
    26181,
    26049,
    25917,
    25785,
    25652,
    25519,
    25385,
    25252,
    25117,
    24983,
    24848,
    24712,
    24576,
    24440,
    24303,
    24166,
    24029,
    23890,
    23752,
    23613,
    23473,
    23333,
    23193,
    23052,
    22910,
    22768,
    22626,
    22482,
    22339,
    22194,
    22049,
    21904,
    21757,
    21611,
    21463,
    21315,
    21166,
    21016,
    20866,
    20715,
    20563,
    20410,
    20257,
    20103,
    19947,
    19791,
    19635,
    19477,
    19318,
    19159,
    18998,
    18836,
    18674,
    18510,
    18345,
    18179,
    18012,
    17844,
    17674,
    17503,
    17331,
    17158,
    16983,
    16807,
    16629,
    16450,
    16269,
    16086,
    15902,
    15716,
    15528,
    15339,
    15147,
    14953,
    14757,
    14559,
    14359,
    14156,
    13951,
    13743,
    13533,
    13319,
    13103,
    12883,
    12660,
    12433,
    12203,
    11969,
    11731,
    11488,
    11240,
    10987,
    10729,
    10466,
    10195,
    9918,
    9634,
    9342,
    9041,
    8730,
    8408,
    8074,
    7727,
    7363,
    6982,
    6579,
    6151,
    5692,
    5194,
    4643,
    4019,
    3280,
    2318,
    0
  };

  //------------------------------------------------------------------------------------------------------
  //
  //------------------------------------------------------------------------------------------------------

  logic [8 : 0] addr0;
  logic [8 : 0] addr1;

  always_ff @(posedge iclk) begin
    if (iclkena) begin
      addr0 <= iaddr0;
      addr1 <= iaddr1;
      //
      odat0 <= cLOG_TAB[addr0];
      odat1 <= cLOG_TAB[addr1];
    end
  end

endmodule
