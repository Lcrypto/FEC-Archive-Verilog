
//
// Project       : ldpc
// Author        : Shekhalev Denis (des00)
// Workfile      : ldpc_parameters.vh
// Description   : LDPC codec parameters and needed functions
//

  //------------------------------------------------------------------------------------------------------
  // Wimax LDPC code parameters matrix parameters
  //------------------------------------------------------------------------------------------------------

  parameter int pCODE   =   5; // coderate = pCODE[3 : 0]/(pCODE[3 : 0]+1), codetype = pCODE[4]
//parameter int pN      = 576;
  parameter int pN      = 2304;

  localparam int pZF    = pN/24 ; // expansion factor

  parameter int pC      = get_H_size(pCODE, 1);
  parameter int pT      = get_H_size(pCODE, 0);

  localparam int cLDPC_NUM  = pT * pZF;
  localparam int cLDPC_DNUM = (pT - pC) * pZF;

  typedef int H_t [pC][pT];

  H_t Hb;

  assign Hb = get_Hb  (pCODE);

  //------------------------------------------------------------------------------------------------------
  // function to get base matrix type
  //------------------------------------------------------------------------------------------------------

  function automatic int get_H_size (input int code, input bit c_nt_sel);
    case (code)
      1 : get_H_size = c_nt_sel ? 12 : 24;
      2 : get_H_size = c_nt_sel ?  8 : 24;
      3 : get_H_size = c_nt_sel ?  6 : 24;
      5 : get_H_size = c_nt_sel ?  4 : 24;
    endcase
  endfunction

  function automatic H_t get_Hb (input int code);
    int Hc_12 [12][24];
    int Hc_23  [8][24];
    int Hc_34  [6][24];
    int Hc_56  [4][24];
    H_t Hc;
  begin
    Hc_12 = '{
              '{-1, 94, 73, -1, -1, -1, -1, -1, 55, 83, -1, -1,  7,  0, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1},
              '{-1, 27, -1, -1, -1, 22, 79,  9, -1, -1, -1, 12, -1,  0,  0, -1, -1, -1, -1, -1, -1, -1, -1, -1},
              '{-1, -1, -1, 24, 22, 81, -1, 33, -1, -1, -1,  0, -1, -1,  0,  0, -1, -1, -1, -1, -1, -1, -1, -1},
              '{61, -1, 47, -1, -1, -1, -1, -1, 65, 25, -1, -1, -1, -1, -1,  0,  0, -1, -1, -1, -1, -1, -1, -1},
              '{-1, -1, 39, -1, -1, -1, 84, -1, -1, 41, 72, -1, -1, -1, -1, -1,  0,  0, -1, -1, -1, -1, -1, -1},
              '{-1, -1, -1, -1, 46, 40, -1, 82, -1, -1, -1, 79,  0, -1, -1, -1, -1,  0,  0, -1, -1, -1, -1, -1},
              '{-1, -1, 95, 53, -1, -1, -1, -1, -1, 14, 18, -1, -1, -1, -1, -1, -1, -1,  0,  0, -1, -1, -1, -1},
              '{-1, 11, 73, -1, -1, -1,  2, -1, -1, 47, -1, -1, -1, -1, -1, -1, -1, -1, -1,  0,  0, -1, -1, -1},
              '{12, -1, -1, -1, 83, 24, -1, 43, -1, -1, -1, 51, -1, -1, -1, -1, -1, -1, -1, -1,  0,  0, -1, -1},
              '{-1, -1, -1, -1, -1, 94, -1, 59, -1, -1, 70, 72, -1, -1, -1, -1, -1, -1, -1, -1, -1,  0,  0, -1},
              '{-1, -1,  7, 65, -1, -1, -1, -1, 39, 49, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1,  0,  0},
              '{43, -1, -1, -1, -1, 66, -1, 41, -1, -1, -1, 26,  7, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1,  0}};

    Hc_23 = '{
              '{ 2, -1, 19, -1, 47, -1, 48, -1, 36, -1, 82, -1, 47, -1, 15, -1, 95,  0, -1, -1, -1, -1, -1, -1},
              '{-1, 69, -1, 88, -1, 33, -1,  3, -1, 16, -1, 37, -1, 40, -1, 48, -1,  0,  0, -1, -1, -1, -1, -1},
              '{10, -1, 86, -1, 62, -1, 28, -1, 85, -1, 16, -1, 34, -1, 73, -1, -1, -1,  0,  0, -1, -1, -1, -1},
              '{-1, 28, -1, 32, -1, 81, -1, 27, -1, 88, -1,  5, -1, 56, -1, 37, -1, -1, -1,  0,  0, -1, -1, -1},
              '{23, -1, 29, -1, 15, -1, 30, -1, 66, -1, 24, -1, 50, -1, 62, -1, -1, -1, -1, -1,  0,  0, -1, -1},
              '{-1, 30, -1, 65, -1, 54, -1, 14, -1,  0, -1, 30, -1, 74, -1,  0, -1, -1, -1, -1, -1,  0,  0, -1},
              '{32, -1,  0, -1, 15, -1, 56, -1, 85, -1,  5, -1,  6, -1, 52, -1,  0, -1, -1, -1, -1, -1,  0,  0},
              '{-1,  0, -1, 47, -1, 13, -1, 61, -1, 84, -1, 55, -1, 78, -1, 41, 95, -1, -1, -1, -1, -1, -1,  0}};

    Hc_34 = '{
              '{ 6, 38,  3, 93, -1, -1, -1, 30, 70, -1, 86, -1, 37, 38,  4, 11, -1, 46, 48,  0, -1, -1, -1, -1},
              '{62, 94, 19, 84, -1, 92, 78, -1, 15, -1, -1, 92, -1, 45, 24, 32, 30, -1, -1,  0,  0, -1, -1, -1},
              '{71, -1, 55, -1, 12, 66, 45, 79, -1, 78, -1, -1, 10, -1, 22, 55, 70, 82, -1, -1,  0,  0, -1, -1},
              '{38, 61, -1, 66,  9, 73, 47, 64, -1, 39, 61, 43, -1, -1, -1, -1, 95, 32,  0, -1, -1,  0,  0, -1},
              '{-1, -1, -1, -1, 32, 52, 55, 80, 95, 22,  6, 51, 24, 90, 44, 20, -1, -1, -1, -1, -1, -1,  0,  0},
              '{-1, 63, 31, 88, 20, -1, -1, -1,  6, 40, 56, 16, 71, 53, -1, -1, 27, 26, 48, -1, -1, -1, -1,  0}};

    Hc_56 = '{
              '{ 1, 25, 55, -1, 47,  4, -1, 91, 84,  8, 86, 52, 82, 33,  5,  0, 36, 20,  4, 77, 80,  0, -1, -1},
              '{-1,  6, -1, 36, 40, 47, 12, 79, 47, -1, 41, 21, 12, 71, 14, 72,  0, 44, 49,  0,  0,  0,  0, -1},
              '{51, 81, 83,  4, 67, -1, 21, -1, 31, 24, 91, 61, 81,  9, 86, 78, 60, 88, 67, 15, -1, -1,  0,  0},
              '{50, -1, 50, 15, -1, 36, 13, 10, 11, 20, 53, 90, 29, 92, 57, 30, 84, 92, 11, 66, 80, -1, -1,  0}};
    //
    for (int j = 0; j < pC; j++) begin
      case (code)
        1 : Hc[j] = Hc_12[j];
        2 : Hc[j] = Hc_23[j];
        3 : Hc[j] = Hc_34[j];
        5 : Hc[j] = Hc_56[j];
      endcase
    end
    //
    for (int i = 0; i < pT; i++) begin
      for (int j = 0; j < pC; j++) begin
        if (Hc[j][i] >= 0)
          get_Hb[j][i] = (Hc[j][i] * pZF)/96;
        else
          get_Hb[j][i] = -1;
      end
    end
    //
//  for (int j = 0; j < pC; j++) begin
//    $display("Hb[%0d] = %p", j, get_Hb[j]);
//  end
  end
  endfunction

