//
// (!!!) IT'S GENERATED FILE for 5/6 coderate, 576 bits do 8 bits per cycle (!!!)
//
  addr_tab[0][0][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[0][0][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[0][0][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[0][1][0] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 127, 127}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[0][1][1] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 127, 127}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[0][1][2] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 2, 2}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[0][2][0] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 127, 127, 127}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[0][2][1] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 2, 2, 2}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[0][2][2] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 127, 127, 127}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[0][3][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][3][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][3][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][4][0] = '{baddr:2, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[0][4][1] = '{baddr:0, offset:'{0, 0, 0, 2, 2, 2, 2, 2}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[0][4][2] = '{baddr:1, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[0][5][0] = '{baddr:1, offset:'{0, 127, 127, 127, 127, 127, 127, 127}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[0][5][1] = '{baddr:2, offset:'{0, 127, 127, 127, 127, 127, 127, 127}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[0][5][2] = '{baddr:0, offset:'{0, 2, 2, 2, 2, 2, 2, 2}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[0][6][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][6][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][6][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][7][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 2, 2}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[0][7][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 127, 127}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[0][7][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 127, 127}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[0][8][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 2, 2, 2}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[0][8][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 127, 127, 127}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[0][8][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 127, 127, 127}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[0][9][0] = '{baddr:1, offset:'{0, 0, 127, 127, 127, 127, 127, 127}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[0][9][1] = '{baddr:2, offset:'{0, 0, 127, 127, 127, 127, 127, 127}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[0][9][2] = '{baddr:0, offset:'{0, 0, 2, 2, 2, 2, 2, 2}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[0][10][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 2, 2, 2}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[0][10][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 127, 127, 127}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[0][10][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 127, 127, 127}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[0][11][0] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 127, 127, 127}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[0][11][1] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 2, 2, 2}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[0][11][2] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 127, 127, 127}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[0][12][0] = '{baddr:0, offset:'{0, 0, 0, 0, 2, 2, 2, 2}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[0][12][1] = '{baddr:1, offset:'{0, 0, 0, 0, 127, 127, 127, 127}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[0][12][2] = '{baddr:2, offset:'{0, 0, 0, 0, 127, 127, 127, 127}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[0][13][0] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[0][13][1] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[0][13][2] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[0][14][0] = '{baddr:1, offset:'{0, 127, 127, 127, 127, 127, 127, 127}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[0][14][1] = '{baddr:2, offset:'{0, 127, 127, 127, 127, 127, 127, 127}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[0][14][2] = '{baddr:0, offset:'{0, 2, 2, 2, 2, 2, 2, 2}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[0][15][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[0][15][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[0][15][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[0][16][0] = '{baddr:2, offset:'{0, 127, 127, 127, 127, 127, 127, 127}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[0][16][1] = '{baddr:0, offset:'{0, 2, 2, 2, 2, 2, 2, 2}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[0][16][2] = '{baddr:1, offset:'{0, 127, 127, 127, 127, 127, 127, 127}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[0][17][0] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 127, 127, 127}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[0][17][1] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 127, 127, 127}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[0][17][2] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 2, 2, 2}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[0][18][0] = '{baddr:1, offset:'{0, 127, 127, 127, 127, 127, 127, 127}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[0][18][1] = '{baddr:2, offset:'{0, 127, 127, 127, 127, 127, 127, 127}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[0][18][2] = '{baddr:0, offset:'{0, 2, 2, 2, 2, 2, 2, 2}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[0][19][0] = '{baddr:0, offset:'{0, 0, 0, 2, 2, 2, 2, 2}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[0][19][1] = '{baddr:1, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[0][19][2] = '{baddr:2, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[0][20][0] = '{baddr:0, offset:'{0, 0, 0, 0, 2, 2, 2, 2}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[0][20][1] = '{baddr:1, offset:'{0, 0, 0, 0, 127, 127, 127, 127}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[0][20][2] = '{baddr:2, offset:'{0, 0, 0, 0, 127, 127, 127, 127}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[0][21][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[0][21][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[0][21][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[0][22][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][22][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][22][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][23][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][23][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[0][23][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[1][0][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[1][0][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[1][0][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[1][1][0] = '{baddr:1, offset:'{0, 127, 127, 127, 127, 127, 127, 127}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[1][1][1] = '{baddr:2, offset:'{0, 127, 127, 127, 127, 127, 127, 127}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[1][1][2] = '{baddr:0, offset:'{0, 2, 2, 2, 2, 2, 2, 2}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[1][2][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[1][2][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[1][2][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[1][3][0] = '{baddr:2, offset:'{0, 127, 127, 127, 127, 127, 127, 127}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[1][3][1] = '{baddr:0, offset:'{0, 2, 2, 2, 2, 2, 2, 2}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[1][3][2] = '{baddr:1, offset:'{0, 127, 127, 127, 127, 127, 127, 127}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[1][4][0] = '{baddr:2, offset:'{0, 0, 127, 127, 127, 127, 127, 127}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[1][4][1] = '{baddr:0, offset:'{0, 0, 2, 2, 2, 2, 2, 2}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[1][4][2] = '{baddr:1, offset:'{0, 0, 127, 127, 127, 127, 127, 127}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[1][5][0] = '{baddr:2, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[1][5][1] = '{baddr:0, offset:'{0, 0, 0, 2, 2, 2, 2, 2}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[1][5][2] = '{baddr:1, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[1][6][0] = '{baddr:1, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[1][6][1] = '{baddr:2, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[1][6][2] = '{baddr:0, offset:'{0, 0, 0, 2, 2, 2, 2, 2}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[1][7][0] = '{baddr:0, offset:'{0, 0, 0, 2, 2, 2, 2, 2}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[1][7][1] = '{baddr:1, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[1][7][2] = '{baddr:2, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[1][8][0] = '{baddr:2, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[1][8][1] = '{baddr:0, offset:'{0, 0, 0, 2, 2, 2, 2, 2}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[1][8][2] = '{baddr:1, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[1][9][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[1][9][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[1][9][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[1][10][0] = '{baddr:2, offset:'{0, 0, 127, 127, 127, 127, 127, 127}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[1][10][1] = '{baddr:0, offset:'{0, 0, 2, 2, 2, 2, 2, 2}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[1][10][2] = '{baddr:1, offset:'{0, 0, 127, 127, 127, 127, 127, 127}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[1][11][0] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 127, 127, 127}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[1][11][1] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 127, 127, 127}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[1][11][2] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 2, 2, 2}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[1][12][0] = '{baddr:1, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[1][12][1] = '{baddr:2, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[1][12][2] = '{baddr:0, offset:'{0, 0, 0, 2, 2, 2, 2, 2}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[1][13][0] = '{baddr:0, offset:'{0, 2, 2, 2, 2, 2, 2, 2}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[1][13][1] = '{baddr:1, offset:'{0, 127, 127, 127, 127, 127, 127, 127}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[1][13][2] = '{baddr:2, offset:'{0, 127, 127, 127, 127, 127, 127, 127}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[1][14][0] = '{baddr:1, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[1][14][1] = '{baddr:2, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[1][14][2] = '{baddr:0, offset:'{0, 0, 0, 2, 2, 2, 2, 2}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[1][15][0] = '{baddr:0, offset:'{0, 0, 2, 2, 2, 2, 2, 2}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[1][15][1] = '{baddr:1, offset:'{0, 0, 127, 127, 127, 127, 127, 127}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[1][15][2] = '{baddr:2, offset:'{0, 0, 127, 127, 127, 127, 127, 127}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[1][16][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][16][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][16][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][17][0] = '{baddr:2, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[1][17][1] = '{baddr:0, offset:'{0, 0, 0, 2, 2, 2, 2, 2}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[1][17][2] = '{baddr:1, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[1][18][0] = '{baddr:2, offset:'{0, 0, 0, 0, 127, 127, 127, 127}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[1][18][1] = '{baddr:0, offset:'{0, 0, 0, 0, 2, 2, 2, 2}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[1][18][2] = '{baddr:1, offset:'{0, 0, 0, 0, 127, 127, 127, 127}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[1][19][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][19][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][19][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][20][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][20][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][20][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][21][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][21][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][21][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][22][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][22][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][22][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[1][23][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[1][23][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[1][23][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][0][0] = '{baddr:2, offset:'{0, 0, 0, 0, 127, 127, 127, 127}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[2][0][1] = '{baddr:0, offset:'{0, 0, 0, 0, 2, 2, 2, 2}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[2][0][2] = '{baddr:1, offset:'{0, 0, 0, 0, 127, 127, 127, 127}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[2][1][0] = '{baddr:0, offset:'{0, 0, 0, 0, 2, 2, 2, 2}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[2][1][1] = '{baddr:1, offset:'{0, 0, 0, 0, 127, 127, 127, 127}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[2][1][2] = '{baddr:2, offset:'{0, 0, 0, 0, 127, 127, 127, 127}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[2][2][0] = '{baddr:0, offset:'{0, 0, 0, 0, 2, 2, 2, 2}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[2][2][1] = '{baddr:1, offset:'{0, 0, 0, 0, 127, 127, 127, 127}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[2][2][2] = '{baddr:2, offset:'{0, 0, 0, 0, 127, 127, 127, 127}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[2][3][0] = '{baddr:1, offset:'{0, 127, 127, 127, 127, 127, 127, 127}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[2][3][1] = '{baddr:2, offset:'{0, 127, 127, 127, 127, 127, 127, 127}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[2][3][2] = '{baddr:0, offset:'{0, 2, 2, 2, 2, 2, 2, 2}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[2][4][0] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[2][4][1] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[2][4][2] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[2][5][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][5][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][5][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][6][0] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 127, 127, 127}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[2][6][1] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 127, 127, 127}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[2][6][2] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 2, 2, 2}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[2][7][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][7][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][7][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][8][0] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][8][1] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][8][2] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][9][0] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 127, 127}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[2][9][1] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 127, 127}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[2][9][2] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 2, 2}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[2][10][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 2, 2}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[2][10][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 127, 127}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[2][10][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 127, 127}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[2][11][0] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][11][1] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][11][2] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][12][0] = '{baddr:0, offset:'{0, 0, 0, 0, 2, 2, 2, 2}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[2][12][1] = '{baddr:1, offset:'{0, 0, 0, 0, 127, 127, 127, 127}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[2][12][2] = '{baddr:2, offset:'{0, 0, 0, 0, 127, 127, 127, 127}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[2][13][0] = '{baddr:1, offset:'{0, 0, 127, 127, 127, 127, 127, 127}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[2][13][1] = '{baddr:2, offset:'{0, 0, 127, 127, 127, 127, 127, 127}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[2][13][2] = '{baddr:0, offset:'{0, 0, 2, 2, 2, 2, 2, 2}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[2][14][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 2, 2, 2}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[2][14][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 127, 127, 127}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[2][14][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 127, 127, 127}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[2][15][0] = '{baddr:0, offset:'{0, 0, 0, 2, 2, 2, 2, 2}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[2][15][1] = '{baddr:1, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[2][15][2] = '{baddr:2, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[2][16][0] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][16][1] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][16][2] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][17][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 2, 2}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[2][17][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 127, 127}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[2][17][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 127, 127}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[2][18][0] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[2][18][1] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[2][18][2] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[2][19][0] = '{baddr:1, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[2][19][1] = '{baddr:2, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[2][19][2] = '{baddr:0, offset:'{0, 0, 0, 2, 2, 2, 2, 2}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[2][20][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][20][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][20][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][21][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][21][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][21][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[2][22][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[2][22][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[2][22][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[2][23][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[2][23][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[2][23][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[3][0][0] = '{baddr:2, offset:'{0, 0, 0, 0, 127, 127, 127, 127}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[3][0][1] = '{baddr:0, offset:'{0, 0, 0, 0, 2, 2, 2, 2}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[3][0][2] = '{baddr:1, offset:'{0, 0, 0, 0, 127, 127, 127, 127}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[3][1][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][1][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][1][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][2][0] = '{baddr:2, offset:'{0, 0, 0, 0, 127, 127, 127, 127}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[3][2][1] = '{baddr:0, offset:'{0, 0, 0, 0, 2, 2, 2, 2}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[3][2][2] = '{baddr:1, offset:'{0, 0, 0, 0, 127, 127, 127, 127}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[3][3][0] = '{baddr:1, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[3][3][1] = '{baddr:2, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[3][3][2] = '{baddr:0, offset:'{0, 0, 0, 2, 2, 2, 2, 2}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[3][4][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][4][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][4][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][5][0] = '{baddr:2, offset:'{0, 127, 127, 127, 127, 127, 127, 127}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[3][5][1] = '{baddr:0, offset:'{0, 2, 2, 2, 2, 2, 2, 2}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[3][5][2] = '{baddr:1, offset:'{0, 127, 127, 127, 127, 127, 127, 127}, sela:'{1, 2, 3, 4, 5, 6, 7, 0}};
  addr_tab[3][6][0] = '{baddr:1, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[3][6][1] = '{baddr:2, offset:'{0, 0, 0, 127, 127, 127, 127, 127}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[3][6][2] = '{baddr:0, offset:'{0, 0, 0, 2, 2, 2, 2, 2}, sela:'{3, 4, 5, 6, 7, 0, 1, 2}};
  addr_tab[3][7][0] = '{baddr:1, offset:'{0, 0, 127, 127, 127, 127, 127, 127}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[3][7][1] = '{baddr:2, offset:'{0, 0, 127, 127, 127, 127, 127, 127}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[3][7][2] = '{baddr:0, offset:'{0, 0, 2, 2, 2, 2, 2, 2}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[3][8][0] = '{baddr:1, offset:'{0, 0, 127, 127, 127, 127, 127, 127}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[3][8][1] = '{baddr:2, offset:'{0, 0, 127, 127, 127, 127, 127, 127}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[3][8][2] = '{baddr:0, offset:'{0, 0, 2, 2, 2, 2, 2, 2}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[3][9][0] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 127, 127, 127}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[3][9][1] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 127, 127, 127}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[3][9][2] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 2, 2, 2}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[3][10][0] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 127, 127, 127}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[3][10][1] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 2, 2, 2}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[3][10][2] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 127, 127, 127}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[3][11][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 2, 2}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[3][11][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 127, 127}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[3][11][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 127, 127}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[3][12][0] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][12][1] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][12][2] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][13][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][13][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][13][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][14][0] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 127, 127}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[3][14][1] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 2, 2}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[3][14][2] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 127, 127}, sela:'{6, 7, 0, 1, 2, 3, 4, 5}};
  addr_tab[3][15][0] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][15][1] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][15][2] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][16][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 2, 2, 2}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[3][16][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 127, 127, 127}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[3][16][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 127, 127, 127}, sela:'{5, 6, 7, 0, 1, 2, 3, 4}};
  addr_tab[3][17][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][17][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][17][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][18][0] = '{baddr:1, offset:'{0, 0, 127, 127, 127, 127, 127, 127}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[3][18][1] = '{baddr:2, offset:'{0, 0, 127, 127, 127, 127, 127, 127}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[3][18][2] = '{baddr:0, offset:'{0, 0, 2, 2, 2, 2, 2, 2}, sela:'{2, 3, 4, 5, 6, 7, 0, 1}};
  addr_tab[3][19][0] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[3][19][1] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[3][19][2] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[3][20][0] = '{baddr:0, offset:'{0, 0, 0, 0, 2, 2, 2, 2}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[3][20][1] = '{baddr:1, offset:'{0, 0, 0, 0, 127, 127, 127, 127}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[3][20][2] = '{baddr:2, offset:'{0, 0, 0, 0, 127, 127, 127, 127}, sela:'{4, 5, 6, 7, 0, 1, 2, 3}};
  addr_tab[3][21][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][21][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][21][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][22][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 2}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][22][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][22][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 127}, sela:'{7, 0, 1, 2, 3, 4, 5, 6}};
  addr_tab[3][23][0] = '{baddr:0, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[3][23][1] = '{baddr:1, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
  addr_tab[3][23][2] = '{baddr:2, offset:'{0, 0, 0, 0, 0, 0, 0, 0}, sela:'{0, 1, 2, 3, 4, 5, 6, 7}};
