/*






  logic          gaus_cordic_tab__iclk       ;
  logic          gaus_cordic_tab__ireset     ;
  logic          gaus_cordic_tab__iclkena    ;
  logic  [8 : 0] gaus_cordic_tab__icos_addr  ;
  logic  [8 : 0] gaus_cordic_tab__isin_addr  ;
  logic [17 : 0] gaus_cordic_tab__ocos       ;
  logic [17 : 0] gaus_cordic_tab__osin       ;



  gaus_cordic_tab
  gaus_cordic_tab
  (
    .iclk      ( gaus_cordic_tab__iclk      ) ,
    .ireset    ( gaus_cordic_tab__ireset    ) ,
    .iclkena   ( gaus_cordic_tab__iclkena   ) ,
    .icos_addr ( gaus_cordic_tab__icos_addr ) ,
    .isin_addr ( gaus_cordic_tab__isin_addr ) ,
    .ocos      ( gaus_cordic_tab__ocos      ) ,
    .osin      ( gaus_cordic_tab__osin      )
  );


  assign gaus_cordic_tab__iclk      = '0 ;
  assign gaus_cordic_tab__ireset    = '0 ;
  assign gaus_cordic_tab__iclkena   = '0 ;
  assign gaus_cordic_tab__icos_addr = '0 ;
  assign gaus_cordic_tab__isin_addr = '0 ;



*/

//
// Project       : gaus_rng
// Author        : Shekhalev Denis (des00)
// Revision      : $Revision$
// Date          : $Date$
// Workfile      : gaus_cordic_tab.v
// Description   : ROM for "cordic"
//

module gaus_cordic_tab
(
  iclk      ,
  ireset    ,
  iclkena   ,
  //
  icos_addr ,
  isin_addr ,
  //
  ocos      ,
  osin
);

  //------------------------------------------------------------------------------------------------------
  //
  //------------------------------------------------------------------------------------------------------

  input  logic          iclk       ;
  input  logic          ireset     ;
  input  logic          iclkena    ;
  //
  input  logic  [8 : 0] icos_addr  ;
  input  logic  [8 : 0] isin_addr  ;
  //
  output logic [17 : 0] ocos       ;
  output logic [17 : 0] osin       ;

  //------------------------------------------------------------------------------------------------------
  //
  //------------------------------------------------------------------------------------------------------

  localparam logic [17 : 0] cCOS_TAB [0 : 511] = '{
    131071,
    131070,
    131066,
    131062,
    131057,
    131050,
    131042,
    131033,
    131022,
    131010,
    130997,
    130983,
    130968,
    130951,
    130933,
    130914,
    130894,
    130872,
    130849,
    130825,
    130800,
    130774,
    130746,
    130717,
    130687,
    130655,
    130623,
    130589,
    130554,
    130517,
    130480,
    130441,
    130401,
    130360,
    130317,
    130273,
    130228,
    130182,
    130135,
    130086,
    130036,
    129985,
    129933,
    129880,
    129825,
    129769,
    129712,
    129653,
    129594,
    129533,
    129471,
    129408,
    129343,
    129277,
    129210,
    129142,
    129073,
    129002,
    128931,
    128858,
    128783,
    128708,
    128631,
    128553,
    128474,
    128394,
    128313,
    128230,
    128146,
    128061,
    127975,
    127887,
    127799,
    127709,
    127617,
    127525,
    127432,
    127337,
    127241,
    127144,
    127046,
    126946,
    126845,
    126744,
    126640,
    126536,
    126431,
    126324,
    126216,
    126107,
    125997,
    125886,
    125773,
    125659,
    125544,
    125428,
    125311,
    125192,
    125073,
    124952,
    124830,
    124706,
    124582,
    124457,
    124330,
    124202,
    124073,
    123943,
    123811,
    123679,
    123545,
    123410,
    123274,
    123137,
    122998,
    122859,
    122718,
    122576,
    122433,
    122289,
    122144,
    121997,
    121850,
    121701,
    121551,
    121400,
    121248,
    121095,
    120940,
    120785,
    120628,
    120470,
    120311,
    120151,
    119990,
    119827,
    119664,
    119499,
    119333,
    119166,
    118998,
    118829,
    118659,
    118488,
    118315,
    118142,
    117967,
    117791,
    117614,
    117436,
    117257,
    117077,
    116895,
    116713,
    116529,
    116345,
    116159,
    115972,
    115784,
    115595,
    115405,
    115214,
    115022,
    114828,
    114634,
    114438,
    114242,
    114044,
    113845,
    113645,
    113445,
    113243,
    113040,
    112836,
    112630,
    112424,
    112217,
    112009,
    111799,
    111589,
    111377,
    111165,
    110951,
    110737,
    110521,
    110304,
    110087,
    109868,
    109648,
    109427,
    109205,
    108982,
    108758,
    108534,
    108308,
    108081,
    107853,
    107624,
    107394,
    107162,
    106930,
    106697,
    106463,
    106228,
    105992,
    105755,
    105517,
    105278,
    105038,
    104797,
    104555,
    104312,
    104068,
    103823,
    103577,
    103330,
    103082,
    102833,
    102584,
    102333,
    102081,
    101828,
    101575,
    101320,
    101064,
    100808,
    100550,
    100292,
    100033,
    99772,
    99511,
    99249,
    98986,
    98722,
    98457,
    98191,
    97924,
    97656,
    97388,
    97118,
    96847,
    96576,
    96304,
    96030,
    95756,
    95481,
    95205,
    94929,
    94651,
    94372,
    94093,
    93812,
    93531,
    93249,
    92966,
    92682,
    92397,
    92111,
    91825,
    91538,
    91249,
    90960,
    90670,
    90379,
    90088,
    89795,
    89502,
    89208,
    88913,
    88617,
    88320,
    88023,
    87724,
    87425,
    87125,
    86824,
    86523,
    86220,
    85917,
    85613,
    85308,
    85002,
    84696,
    84388,
    84080,
    83771,
    83462,
    83151,
    82840,
    82528,
    82215,
    81902,
    81587,
    81272,
    80956,
    80640,
    80322,
    80004,
    79685,
    79366,
    79045,
    78724,
    78402,
    78079,
    77756,
    77432,
    77107,
    76782,
    76455,
    76128,
    75801,
    75472,
    75143,
    74813,
    74483,
    74152,
    73820,
    73487,
    73154,
    72820,
    72485,
    72150,
    71814,
    71477,
    71139,
    70801,
    70463,
    70123,
    69783,
    69442,
    69101,
    68759,
    68416,
    68073,
    67729,
    67384,
    67039,
    66693,
    66347,
    66000,
    65652,
    65304,
    64955,
    64605,
    64255,
    63904,
    63553,
    63201,
    62848,
    62495,
    62141,
    61787,
    61432,
    61076,
    60720,
    60364,
    60007,
    59649,
    59290,
    58931,
    58572,
    58212,
    57851,
    57490,
    57129,
    56766,
    56404,
    56041,
    55677,
    55312,
    54948,
    54582,
    54216,
    53850,
    53483,
    53116,
    52748,
    52380,
    52011,
    51641,
    51271,
    50901,
    50530,
    50159,
    49787,
    49415,
    49042,
    48669,
    48296,
    47922,
    47547,
    47172,
    46797,
    46421,
    46045,
    45668,
    45291,
    44913,
    44535,
    44157,
    43778,
    43399,
    43019,
    42639,
    42259,
    41878,
    41497,
    41115,
    40733,
    40350,
    39968,
    39585,
    39201,
    38817,
    38433,
    38048,
    37663,
    37278,
    36892,
    36506,
    36120,
    35733,
    35346,
    34959,
    34571,
    34183,
    33794,
    33406,
    33017,
    32627,
    32238,
    31848,
    31458,
    31067,
    30676,
    30285,
    29894,
    29502,
    29110,
    28718,
    28326,
    27933,
    27540,
    27147,
    26753,
    26359,
    25965,
    25571,
    25176,
    24782,
    24387,
    23991,
    23596,
    23200,
    22804,
    22408,
    22012,
    21615,
    21219,
    20822,
    20425,
    20027,
    19630,
    19232,
    18834,
    18436,
    18038,
    17640,
    17241,
    16843,
    16444,
    16045,
    15645,
    15246,
    14847,
    14447,
    14047,
    13647,
    13247,
    12847,
    12447,
    12047,
    11646,
    11246,
    10845,
    10444,
    10043,
    9642,
    9241,
    8840,
    8439,
    8037,
    7636,
    7235,
    6833,
    6431,
    6030,
    5628,
    5226,
    4824,
    4423,
    4021,
    3619,
    3217,
    2815,
    2413,
    2011,
    1608,
    1206,
    804,
    402,
    0
  };

  //------------------------------------------------------------------------------------------------------
  //
  //------------------------------------------------------------------------------------------------------

  logic [10 : 0] cos_addr  ;
  logic [10 : 0] sin_addr  ;

  always_ff @(posedge iclk) begin
    if (iclkena) begin
      cos_addr <= icos_addr;
      sin_addr <= isin_addr;
      //
      ocos     <= cCOS_TAB[cos_addr];
      osin     <= cCOS_TAB[sin_addr];
    end
  end

endmodule
