//
// Project       : bch
// Author        : Shekhalev Denis (des00)
// Revision      : $Revision: 12476 $
// Date          : $Date$
// Workfile      : rs_define.vh
// Description   : rs modules macros file
//

//`define __RS_BERLEKAMP_DEBUG_LOG__
//`define __RS_CHIENY_DEBUG_LOG__
